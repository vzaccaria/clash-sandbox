-- Automatically generated VHDL
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use work.all;
use work.types.all;

entity shift1_5 is
  port(i_i1     : in array_of_unsigned_8(0 to 15);
       topLet_o : out array_of_unsigned_8(0 to 15));
end;

architecture structural of shift1_5 is
  signal repANF_0  : unsigned(7 downto 0);
  signal repANF_1  : unsigned(7 downto 0);
  signal repANF_2  : unsigned(7 downto 0);
  signal repANF_3  : unsigned(7 downto 0);
  signal repANF_4  : unsigned(7 downto 0);
  signal repANF_5  : unsigned(7 downto 0);
  signal repANF_6  : unsigned(7 downto 0);
  signal repANF_7  : unsigned(7 downto 0);
  signal repANF_8  : unsigned(7 downto 0);
  signal repANF_9  : unsigned(7 downto 0);
  signal repANF_10 : unsigned(7 downto 0);
  signal repANF_11 : unsigned(7 downto 0);
  signal repANF_12 : unsigned(7 downto 0);
  signal repANF_13 : unsigned(7 downto 0);
  signal repANF_14 : unsigned(7 downto 0);
  signal repANF_15 : unsigned(7 downto 0);
  signal repANF_16 : array_of_unsigned_8(0 to 0);
  signal repANF_17 : array_of_unsigned_8(0 to 1);
  signal repANF_18 : array_of_unsigned_8(0 to 2);
  signal repANF_19 : array_of_unsigned_8(0 to 3);
  signal repANF_20 : array_of_unsigned_8(0 to 4);
  signal repANF_21 : array_of_unsigned_8(0 to 5);
  signal repANF_22 : array_of_unsigned_8(0 to 6);
  signal repANF_23 : array_of_unsigned_8(0 to 7);
  signal repANF_24 : array_of_unsigned_8(0 to 8);
  signal repANF_25 : array_of_unsigned_8(0 to 9);
  signal repANF_26 : array_of_unsigned_8(0 to 10);
  signal repANF_27 : array_of_unsigned_8(0 to 11);
  signal repANF_28 : array_of_unsigned_8(0 to 12);
  signal repANF_29 : array_of_unsigned_8(0 to 13);
  signal repANF_30 : array_of_unsigned_8(0 to 14);
  signal tmp_31    : unsigned(7 downto 0);
  signal tmp_35    : unsigned(7 downto 0);
  signal tmp_39    : unsigned(7 downto 0);
  signal tmp_43    : unsigned(7 downto 0);
  signal tmp_47    : unsigned(7 downto 0);
  signal tmp_51    : unsigned(7 downto 0);
  signal tmp_55    : unsigned(7 downto 0);
  signal tmp_59    : unsigned(7 downto 0);
  signal tmp_63    : unsigned(7 downto 0);
  signal tmp_67    : unsigned(7 downto 0);
  signal tmp_71    : unsigned(7 downto 0);
  signal tmp_75    : unsigned(7 downto 0);
  signal tmp_79    : unsigned(7 downto 0);
  signal tmp_83    : unsigned(7 downto 0);
  signal tmp_87    : unsigned(7 downto 0);
  signal tmp_91    : unsigned(7 downto 0);
begin
  indexVec_n_32 : block
    signal n_33 : array_of_unsigned_8(0 to 15);
    signal n_34 : integer;
  begin
    n_33 <= i_i1;
    n_34 <= 0;
    -- pragma translate_off
    process (n_33,n_34)
    begin
      if n_34 < n_33'low or n_34 > n_33'high then
        assert false report ("Index: " & integer'image(n_34) & ", is out of bounds: " & integer'image(n_33'low) & " to " & integer'image(n_33'high)) severity warning;
        tmp_31 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_31 <= n_33(n_34);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_0 <= tmp_31;
  
  indexVec_n_36 : block
    signal n_37 : array_of_unsigned_8(0 to 15);
    signal n_38 : integer;
  begin
    n_37 <= i_i1;
    n_38 <= 5;
    -- pragma translate_off
    process (n_37,n_38)
    begin
      if n_38 < n_37'low or n_38 > n_37'high then
        assert false report ("Index: " & integer'image(n_38) & ", is out of bounds: " & integer'image(n_37'low) & " to " & integer'image(n_37'high)) severity warning;
        tmp_35 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_35 <= n_37(n_38);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_1 <= tmp_35;
  
  indexVec_n_40 : block
    signal n_41 : array_of_unsigned_8(0 to 15);
    signal n_42 : integer;
  begin
    n_41 <= i_i1;
    n_42 <= 10;
    -- pragma translate_off
    process (n_41,n_42)
    begin
      if n_42 < n_41'low or n_42 > n_41'high then
        assert false report ("Index: " & integer'image(n_42) & ", is out of bounds: " & integer'image(n_41'low) & " to " & integer'image(n_41'high)) severity warning;
        tmp_39 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_39 <= n_41(n_42);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_2 <= tmp_39;
  
  indexVec_n_44 : block
    signal n_45 : array_of_unsigned_8(0 to 15);
    signal n_46 : integer;
  begin
    n_45 <= i_i1;
    n_46 <= 15;
    -- pragma translate_off
    process (n_45,n_46)
    begin
      if n_46 < n_45'low or n_46 > n_45'high then
        assert false report ("Index: " & integer'image(n_46) & ", is out of bounds: " & integer'image(n_45'low) & " to " & integer'image(n_45'high)) severity warning;
        tmp_43 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_43 <= n_45(n_46);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_3 <= tmp_43;
  
  indexVec_n_48 : block
    signal n_49 : array_of_unsigned_8(0 to 15);
    signal n_50 : integer;
  begin
    n_49 <= i_i1;
    n_50 <= 4;
    -- pragma translate_off
    process (n_49,n_50)
    begin
      if n_50 < n_49'low or n_50 > n_49'high then
        assert false report ("Index: " & integer'image(n_50) & ", is out of bounds: " & integer'image(n_49'low) & " to " & integer'image(n_49'high)) severity warning;
        tmp_47 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_47 <= n_49(n_50);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_4 <= tmp_47;
  
  indexVec_n_52 : block
    signal n_53 : array_of_unsigned_8(0 to 15);
    signal n_54 : integer;
  begin
    n_53 <= i_i1;
    n_54 <= 9;
    -- pragma translate_off
    process (n_53,n_54)
    begin
      if n_54 < n_53'low or n_54 > n_53'high then
        assert false report ("Index: " & integer'image(n_54) & ", is out of bounds: " & integer'image(n_53'low) & " to " & integer'image(n_53'high)) severity warning;
        tmp_51 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_51 <= n_53(n_54);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_5 <= tmp_51;
  
  indexVec_n_56 : block
    signal n_57 : array_of_unsigned_8(0 to 15);
    signal n_58 : integer;
  begin
    n_57 <= i_i1;
    n_58 <= 14;
    -- pragma translate_off
    process (n_57,n_58)
    begin
      if n_58 < n_57'low or n_58 > n_57'high then
        assert false report ("Index: " & integer'image(n_58) & ", is out of bounds: " & integer'image(n_57'low) & " to " & integer'image(n_57'high)) severity warning;
        tmp_55 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_55 <= n_57(n_58);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_6 <= tmp_55;
  
  indexVec_n_60 : block
    signal n_61 : array_of_unsigned_8(0 to 15);
    signal n_62 : integer;
  begin
    n_61 <= i_i1;
    n_62 <= 3;
    -- pragma translate_off
    process (n_61,n_62)
    begin
      if n_62 < n_61'low or n_62 > n_61'high then
        assert false report ("Index: " & integer'image(n_62) & ", is out of bounds: " & integer'image(n_61'low) & " to " & integer'image(n_61'high)) severity warning;
        tmp_59 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_59 <= n_61(n_62);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_7 <= tmp_59;
  
  indexVec_n_64 : block
    signal n_65 : array_of_unsigned_8(0 to 15);
    signal n_66 : integer;
  begin
    n_65 <= i_i1;
    n_66 <= 8;
    -- pragma translate_off
    process (n_65,n_66)
    begin
      if n_66 < n_65'low or n_66 > n_65'high then
        assert false report ("Index: " & integer'image(n_66) & ", is out of bounds: " & integer'image(n_65'low) & " to " & integer'image(n_65'high)) severity warning;
        tmp_63 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_63 <= n_65(n_66);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_8 <= tmp_63;
  
  indexVec_n_68 : block
    signal n_69 : array_of_unsigned_8(0 to 15);
    signal n_70 : integer;
  begin
    n_69 <= i_i1;
    n_70 <= 13;
    -- pragma translate_off
    process (n_69,n_70)
    begin
      if n_70 < n_69'low or n_70 > n_69'high then
        assert false report ("Index: " & integer'image(n_70) & ", is out of bounds: " & integer'image(n_69'low) & " to " & integer'image(n_69'high)) severity warning;
        tmp_67 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_67 <= n_69(n_70);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_9 <= tmp_67;
  
  indexVec_n_72 : block
    signal n_73 : array_of_unsigned_8(0 to 15);
    signal n_74 : integer;
  begin
    n_73 <= i_i1;
    n_74 <= 2;
    -- pragma translate_off
    process (n_73,n_74)
    begin
      if n_74 < n_73'low or n_74 > n_73'high then
        assert false report ("Index: " & integer'image(n_74) & ", is out of bounds: " & integer'image(n_73'low) & " to " & integer'image(n_73'high)) severity warning;
        tmp_71 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_71 <= n_73(n_74);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_10 <= tmp_71;
  
  indexVec_n_76 : block
    signal n_77 : array_of_unsigned_8(0 to 15);
    signal n_78 : integer;
  begin
    n_77 <= i_i1;
    n_78 <= 7;
    -- pragma translate_off
    process (n_77,n_78)
    begin
      if n_78 < n_77'low or n_78 > n_77'high then
        assert false report ("Index: " & integer'image(n_78) & ", is out of bounds: " & integer'image(n_77'low) & " to " & integer'image(n_77'high)) severity warning;
        tmp_75 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_75 <= n_77(n_78);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_11 <= tmp_75;
  
  indexVec_n_80 : block
    signal n_81 : array_of_unsigned_8(0 to 15);
    signal n_82 : integer;
  begin
    n_81 <= i_i1;
    n_82 <= 12;
    -- pragma translate_off
    process (n_81,n_82)
    begin
      if n_82 < n_81'low or n_82 > n_81'high then
        assert false report ("Index: " & integer'image(n_82) & ", is out of bounds: " & integer'image(n_81'low) & " to " & integer'image(n_81'high)) severity warning;
        tmp_79 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_79 <= n_81(n_82);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_12 <= tmp_79;
  
  indexVec_n_84 : block
    signal n_85 : array_of_unsigned_8(0 to 15);
    signal n_86 : integer;
  begin
    n_85 <= i_i1;
    n_86 <= 1;
    -- pragma translate_off
    process (n_85,n_86)
    begin
      if n_86 < n_85'low or n_86 > n_85'high then
        assert false report ("Index: " & integer'image(n_86) & ", is out of bounds: " & integer'image(n_85'low) & " to " & integer'image(n_85'high)) severity warning;
        tmp_83 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_83 <= n_85(n_86);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_13 <= tmp_83;
  
  indexVec_n_88 : block
    signal n_89 : array_of_unsigned_8(0 to 15);
    signal n_90 : integer;
  begin
    n_89 <= i_i1;
    n_90 <= 6;
    -- pragma translate_off
    process (n_89,n_90)
    begin
      if n_90 < n_89'low or n_90 > n_89'high then
        assert false report ("Index: " & integer'image(n_90) & ", is out of bounds: " & integer'image(n_89'low) & " to " & integer'image(n_89'high)) severity warning;
        tmp_87 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_87 <= n_89(n_90);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_14 <= tmp_87;
  
  indexVec_n_92 : block
    signal n_93 : array_of_unsigned_8(0 to 15);
    signal n_94 : integer;
  begin
    n_93 <= i_i1;
    n_94 <= 11;
    -- pragma translate_off
    process (n_93,n_94)
    begin
      if n_94 < n_93'low or n_94 > n_93'high then
        assert false report ("Index: " & integer'image(n_94) & ", is out of bounds: " & integer'image(n_93'low) & " to " & integer'image(n_93'high)) severity warning;
        tmp_91 <= (others => 'X');
      else
      -- pragma translate_on
        tmp_91 <= n_93(n_94);
      -- pragma translate_off
      end if;
    end process;
    -- pragma translate_on
  end block;
  
  repANF_15 <= tmp_91;
  
  repANF_16 <= array_of_unsigned_8'(0 => repANF_15);
  
  repANF_17 <= array_of_unsigned_8'(unsigned'(repANF_14) & repANF_16);
  
  repANF_18 <= array_of_unsigned_8'(unsigned'(repANF_13) & repANF_17);
  
  repANF_19 <= array_of_unsigned_8'(unsigned'(repANF_12) & repANF_18);
  
  repANF_20 <= array_of_unsigned_8'(unsigned'(repANF_11) & repANF_19);
  
  repANF_21 <= array_of_unsigned_8'(unsigned'(repANF_10) & repANF_20);
  
  repANF_22 <= array_of_unsigned_8'(unsigned'(repANF_9) & repANF_21);
  
  repANF_23 <= array_of_unsigned_8'(unsigned'(repANF_8) & repANF_22);
  
  repANF_24 <= array_of_unsigned_8'(unsigned'(repANF_7) & repANF_23);
  
  repANF_25 <= array_of_unsigned_8'(unsigned'(repANF_6) & repANF_24);
  
  repANF_26 <= array_of_unsigned_8'(unsigned'(repANF_5) & repANF_25);
  
  repANF_27 <= array_of_unsigned_8'(unsigned'(repANF_4) & repANF_26);
  
  repANF_28 <= array_of_unsigned_8'(unsigned'(repANF_3) & repANF_27);
  
  repANF_29 <= array_of_unsigned_8'(unsigned'(repANF_2) & repANF_28);
  
  repANF_30 <= array_of_unsigned_8'(unsigned'(repANF_1) & repANF_29);
  
  topLet_o <= array_of_unsigned_8'(unsigned'(repANF_0) & repANF_30);
end;
